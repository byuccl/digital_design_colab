module StateMachine(
  //Signals
);
  
endmodule
