module circuit(

);


endmodule
